`timescale 1ns/1ps

`include "../../include/global.svh"

module dcache(
);
    
endmodule